`define MM_RAM_DEPTH 64
`define CONST0_RAM_DEPTH 64
`define CONST1_RAM_DEPTH 64
`define ADD0_RAM_DEPTH 64
`define ADD1_RAM_DEPTH 64
`define ADD2_RAM_DEPTH 64
`define ADD3_RAM_DEPTH 64
`define ADD4_RAM_DEPTH 64
`define ADD5_RAM_DEPTH 64
`define ADD6_RAM_DEPTH 64
`define ADD7_RAM_DEPTH 64

`define MM_RAM_SIZE 6
`define CONST0_RAM_SIZE 6
`define CONST1_RAM_SIZE 6
`define ADD0_RAM_SIZE 6
`define ADD1_RAM_SIZE 6
`define ADD2_RAM_SIZE 6
`define ADD3_RAM_SIZE 6
`define ADD4_RAM_SIZE 6
`define ADD5_RAM_SIZE 6
`define ADD6_RAM_SIZE 6
`define ADD7_RAM_SIZE 6

`define OPR_NUM_SIZE    4  // log(10)
`define MM0     0
`define CONST0  1
`define CONST1  2
`define ADD0    3
`define ADD1    4
`define ADD2    5
`define ADD3    6
`define ADD4    7
`define ADD5    8
`define ADD6    9
`define ADD7    10
`define CALC_STATE_SIZE 7
`define CALC_CONJ_STATE_SIZE `CALC_STATE_SIZE'd4
`define CALC_FROB_STATE_SIZE `CALC_STATE_SIZE'd16
`define CALC_INV_STATE_SIZE `CALC_STATE_SIZE'd106
`define CALC_MUL_STATE_SIZE `CALC_STATE_SIZE'd34
`define CALC_MUL_CONJ_STATE_SIZE `CALC_STATE_SIZE'd34
`define CALC_PADD_STATE_SIZE `CALC_STATE_SIZE'd46
`define CALC_PDBL_STATE_SIZE `CALC_STATE_SIZE'd36
`define CALC_PMINUS_STATE_SIZE `CALC_STATE_SIZE'd46
`define CALC_SPARSE_STATE_SIZE `CALC_STATE_SIZE'd25
`define CALC_SQR_STATE_SIZE `CALC_STATE_SIZE'd26
`define CALC_SQR012345_STATE_SIZE `CALC_STATE_SIZE'd20
